
-- 32 BIT MEMORY

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;



------------------------------- ENTITIY -------------------------------------------

ENTITY insmem IS
    PORT(din : IN std_logic_vector(31 DOWNTO 0);
         addr: IN std_logic_vector(31 DOWNTO 0);
         nrw : IN std_logic;
         dout: OUT std_logic_vector(31 DOWNTO 0)
         );
END insmem;


------------------------------- ARCHITECTURE ------------------------------------------


ARCHITECTURE mem OF insmem IS

    TYPE reg_bank IS ARRAY (0 TO 31) OF std_logic_vector(31 DOWNTO 0);
    SIGNAL buff : reg_bank;
    
BEGIN

    PROCESS (addr,din,nrw)
    BEGIN
        IF nrw='0' THEN
            dout<=buff(conv_integer(addr));
            buff(0)  <= "00000000000000000000100000100100" ;
            buff(1)  <= "00000000000000000000100000100100" ;
            buff(2)  <= "00000000000000000001000000100100" ;
            buff(3)  <= "00000000001000100001100000100001" ;
            buff(4)  <= "00000000010000110010000000100110" ;
            buff(5)  <= "00000000000000010010100000101011" ;
            buff(6)  <= "00000000000000010011000011000010" ;
            buff(7)  <= "00000000000000110011100000000110" ;
            buff(8)  <= "00000000000001000100000000100011" ;
            buff(9)  <= "00000000000000110100100000100101" ;
            buff(10) <= "00000000000001110101001100000000" ;
            buff(11) <= "00000000111010000101100000000100" ;
            buff(12) <= "00000000000000000110000000100100" ;
            buff(13) <= "00000000001000100110100000100001" ;
            buff(14) <= "00000000010000110111000000100110" ;
            buff(15) <= "00000000000000010111100000101011" ;
            buff(16) <= "00000000000000011000000011000010" ;
            buff(17) <= "00000000000000111000100000000110" ;
            buff(18) <= "00000000000001001001000000100011" ;
            buff(19) <= "00000000000000111001100000100101" ;
            buff(20) <= "00000000000001111010001100000000" ;
            buff(21) <= "00000000111010001010100000000100" ;
            buff(22) <= "00000000000000001011000000100100" ;
            buff(23) <= "00000000001000101011100000100001" ;
            buff(24) <= "00000000010000111100000000100110" ;
            buff(25) <= "00000000000000011100100000101011" ;
            buff(26) <= "00000000000000011101000011000010" ;
            buff(27) <= "00000000000000111101100000000110" ;
            buff(28) <= "00000000000001001110000000100011" ;
            buff(29) <= "00000000000000111110100000100101" ;
            buff(30) <= "00000000000001111111001100000000" ;
            buff(31) <= "00000000111010001111100000000100" ;
        ELSE
            buff(conv_integer(addr))<=din;
        END IF;
    END PROCESS;
END mem;







